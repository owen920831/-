`timescale 1ns/1ps

module Majority(a, b, c, out);
input a, b, c;
output out;

endmodule